module hex_7s (
	input  [3:0] H,
	output reg [6:0] S);
	always@(H)
	case (H)  //ANODO COMUN
		0:  S = 7'b0000001;
		1:  S = 7'b1001111;
		2:  S = 7'b0010010;
		3:  S = 7'b0000110;
		4:  S = 7'b1001100;
		5:  S = 7'b0100100;
		6:  S = 7'b0100000;
		7:  S = 7'b0001111;
		8:  S = 7'b0000000;
		9:  S = 7'b0001100;
		10: S = 7'b0001000;
		11: S = 7'b1100000;
		12: S = 7'b0110001;
		13: S = 7'b1000010;
		14: S = 7'b0110000;
		15: S = 7'b0111000;
	endcase
endmodule
